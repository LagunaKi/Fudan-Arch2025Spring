`ifndef __FETCH_SV
`define __FETHC_SV

`ifdef VERILATOR
`include "include/common.sv"
`include "include/pipes.sv"
`else

`endif 

module fetch 
    import common::*;
    import pipes::*;(

    output fetch_data_t dataF, // fetch_data_t defined in pipes.sv
    input u32 raw_instr
);

    assign dataF.raw_instr = raw_instr;

endmodule



`endif


