`ifndef __CORE_SV
`define __CORE_SV

`ifdef VERILATOR
`include "include/csr.sv"
`include "include/common.sv"
`include "pipeline/fetch/fetch.sv"
`include "pipeline/fetch/pcselect.sv"
`include "pipeline/decode/decode.sv"
`include "pipeline/execute/execute.sv"
`include "pipeline/memory/memory.sv"
`include "pipeline/memory/mmu.sv"
`include "pipeline/writeback/writeback.sv"
`include "pipeline/regfile/regfile.sv"
`include "pipeline/regfile/csr_regfile.sv"
`include "pipeline/regs/reg_FD.sv"
`include "pipeline/regs/reg_DE.sv"
`include "pipeline/regs/reg_EM.sv"
`include "pipeline/regs/reg_MW.sv"

`endif

module core 
	import csr_pkg::*;
	import common::*;
(
	input logic clk, reset,
	output ibus_req_t  ireq,
	input  ibus_resp_t iresp,
	output dbus_req_t  dreq,
	input  dbus_resp_t dresp,
	input logic trint, swint, exint
);

    /* TODO: Add your CPU-Core here. */

    u64       pc, pc_nxt, offset;
    u32       raw_instr;
    u1        handin;
    fetch_data_t       dataF, dataF_nxt, saved_dataF;
    decode_data_t      dataD, dataD_nxt;
    execute_data_t     dataE, dataE_nxt;
    memory_data_t      dataM, dataM_nxt;
    writeback_data_t   dataW;
    creg_addr_t        ra1, ra2;
    word_t             rd1, rd2, csr_rd;
	csr_addr_t         csr_ra;
    u1                 stallpc, stalldata, stall, bubble, flush, csr_write;
	u1 				   hazard_ra1, hazard_ra2, hazard_jalr, hazard_csr;
	instfunc_t         op_in, op_out;
    
    // MMU signals
    u1 mmu_page_fault;
    dbus_req_t mmu_dreq;
    ibus_req_t mmu_ireq;
    dbus_resp_t mmu_dresp;
    ibus_resp_t mmu_iresp;

    u2 privilege_mode;
    u2 privilege_mode_nxt;

    assign stallpc = mmu_ireq.valid & (~mmu_iresp.data_ok);
	assign stalldata = mmu_dreq.valid & (~mmu_dresp.data_ok);
	assign stall = dataD.stall;
	assign handin = ~dataW.stall;

    always_ff @(posedge clk) begin
        if (reset) begin
            pc <= 64'h8000_0000;
            // mmu_ireq.addr <= '0;
            mmu_ireq.addr <= 64'h8000_0000;
            mmu_ireq.valid <= '1;
        end 
		else begin
            pc <= pc_nxt;
            if (mmu_ireq.valid == 1'b0) begin
                mmu_ireq.addr <= pc_nxt;
                mmu_ireq.valid <= 1'b1;
            end 
			else begin
                if (mmu_iresp.data_ok == 0) begin
                    mmu_ireq.addr <= mmu_ireq.addr;
                    mmu_ireq.valid <= mmu_ireq.valid;
                end 
				else begin
                    mmu_ireq.addr <= mmu_ireq.addr;
                    mmu_ireq.valid <= 1'b0;
                end
            end
        end
    end

	always_comb begin
		if(bubble)begin
			raw_instr = '0;
		end
		else begin
        	raw_instr = (mmu_iresp.data_ok == 1) ? mmu_iresp.data : '0;
		end
    end

	// Pipeline flush control
    assign csr_write = (dataW.ctl.op inside {CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI, ECALL, MRET}) & ~dataW.stall;
    
    assign flush = csr_write;

	// data hazard
    // CSR hazard detection
    assign hazard_csr = (~stall) && (
        (dataD.ctl.op inside {CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI}) &&
        ((~dataE.stall && dataE.ctl.op inside {CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI} && 
          dataD.ctl.csr_ops[0].addr == dataE.ctl.csr_ops[0].addr) ||
         (~dataM.stall && dataM.ctl.op inside {CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI} &&
          dataD.ctl.csr_ops[0].addr == dataM.ctl.csr_ops[0].addr) ||
         (~dataW.stall && dataW.ctl.op inside {CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI} &&
          dataD.ctl.csr_ops[0].addr == dataW.ctl.csr_ops[0].addr))
    );

	assign hazard_ra1 = (~stall) && (
						(~dataE.stall && ra1 == dataE.dst) || 
						(~dataM.stall && ra1 == dataM.dst) || 
						(~dataW.stall && ra1 == dataW.dst));

	assign hazard_ra2 = (~stall) && (
						(~dataE.stall && ra2 == dataE.dst) || 
						(~dataM.stall && ra2 == dataM.dst) || 
						(~dataW.stall && ra2 == dataW.dst));
	
	assign hazard_jalr = (~stall && dataD.ctl.op == JALR) && (
						(~dataE.stall && ra1 == dataE.dst) ||
						(~dataM.stall && ra1 == dataM.dst) ||
						(~dataW.stall && ra1 == dataW.dst));

	assign bubble = hazard_ra1 || hazard_ra2 || hazard_jalr || hazard_csr;
	// assign bubble = hazard_ra1 || hazard_ra2;

	always_comb begin
		if(dataD.ctl.op == JALR)begin
			if(hazard_jalr)begin
				op_out = MAINTAIN;
			end
			else begin
				op_out = F_JALR;
			end
		end
		else begin
			op_out = op_in;
		end
	end


    pcselect pcselect (
		.pc, .stalldata, .stallpc, 
        //.ireq,
        .ireq(mmu_ireq),
		.pc_selected(pc_nxt),
		.stall, .bubble, .flush, 
		.op(op_out), .offset,
		.mepc(csr_regfile.mepc_nxt),  // Connect MEPC from CSR
        .mtvec(csr_regfile.mtvec_nxt) // Connect MTVEC from CSR
	);


    fetch fetch (
        .raw_instr, 
        // .ireq,
        .ireq(mmu_ireq), 
        .pc, .dataF
    );

    reg_FD reg_FD (
        .clk,  .reset , .ireq, .flush, 
		.stallpc, .stalldata,
		.saved_dataF_in (saved_dataF),
		.saved_dataF_out (saved_dataF), 
		.last_dataF (dataF_nxt),
        .dataF_in       (dataF),
        .dataF_out      (dataF_nxt),
		.bubble
    );

    decode decode (
        .dataF  (dataF_nxt),
        .dataD,
        .ra1, .ra2,
        .rd1, .rd2, .csr_rd, 
		.op     (op_in),
		.offset, .csr_ra
    );

    reg_DE reg_DE (
        .clk ,.reset , .stalldata, .flush, 
        .dataD_in   (dataD),
        .dataD_out  (dataD_nxt),
		.last_dataD (dataD_nxt),
		.bubble
    );

    execute execute (
        .clk            (clk),
        .reset          (reset),
        .dataD          (dataD_nxt),
        .dataE          (dataE),
        .privilege_mode (privilege_mode)
    );

    reg_EM reg_EM (
        .clk, .reset, .stalldata, .flush, 
        .dataE_in       (dataE),
        .dataE_out      (dataE_nxt),
		.last_dataE     (dataE_nxt)
    );

    always_comb begin
        privilege_mode_nxt = privilege_mode;
        if(reset)begin
            privilege_mode_nxt = PRIVILEGE_M_MODE;
        end
        else if(dataW.ctl.is_mret & ~stallpc)begin //prevent m_mode ireq handled in u_mode
            privilege_mode_nxt = (csr_regfile.mstatus_nxt[12:11] == 2'b11) ? PRIVILEGE_M_MODE :
                                (csr_regfile.mstatus_nxt[12:11] == 2'b01) ? PRIVILEGE_S_MODE :
                                PRIVILEGE_U_MODE;
        end
        else if(dataW.ctl.is_ecall)begin
            privilege_mode_nxt = PRIVILEGE_M_MODE;
        end
    end

    always_ff @(posedge clk) begin
        if (reset) begin
            privilege_mode <= PRIVILEGE_M_MODE;
        end 
		else begin
            privilege_mode <= privilege_mode_nxt;
        end
    end

    mmu mmu (
        .clk            (clk),
        .reset          (reset),
        .privilege_mode (privilege_mode),
        .satp           (csr_regfile.satp_nxt),
        .dreq           (dreq),
        .mmu_dreq       (mmu_dreq),
        .ireq           (ireq),
        .mmu_ireq       (mmu_ireq),
        .mmu_page_fault (mmu_page_fault),
        .dresp          (dresp),
        .iresp          (iresp),
        .mmu_dresp      (mmu_dresp),
        .mmu_iresp      (mmu_iresp)
    );

    memory memory(
        .dataE(dataE_nxt),               // Unchanged pipeline data
        .dresp(mmu_dresp), // Responses go through MMU
        // .dreq(dreq),                    // Memory requests go directly to system
        .dreq(mmu_dreq),
        .dataM(dataM),                  // Unchanged pipeline output
        .mmu_page_fault(mmu_page_fault) // MMU page fault signal
    );

    // always_comb begin
    //     // Default assignments
    //     dataM.exception = 1'b0;
    //     dataM.cause = '0;
    //     dataM.tval = '0;
        
    //     if (mmu_page_fault) begin
    //         dataM.exception = 1'b1;
    //         dataM.cause = dataE_nxt.ctl.memwrite ? STORE_PAGE_FAULT : LOAD_PAGE_FAULT;
    //         dataM.tval = dataE_nxt.mem_addr;
    //     end
    // end

    reg_MW reg_MW (
        .clk, .reset, .stalldata, .flush, 
        .dataM_in       (dataM),
        .dataM_out      (dataM_nxt),
		.last_dataM (dataM_nxt)
    );

    writeback writeback (
        .dataM          (dataM_nxt),
        .dataW          (dataW)
    );

    // CSR register file
    csr_regfile csr_regfile (
        .clk            (clk),
        .reset          (reset),
        // Multi-register write port (for MRET/ECALL)
        .csr_ops     (dataW.ctl.csr_ops),
        // Read port
        .ra          (csr_ra),
        .rd          (csr_rd)
    );

    regfile regfile (
        .clk            (clk),
        .reset          (reset),
        .ra1            (ra1),
        .ra2            (ra2),
        .rd1            (rd1),
        .rd2            (rd2),
        .WE             (dataW.ctl.regwrite & ~dataW.stall),
        .wa             (dataW.dst),
        .wd             (dataW.result)
    );


    


`ifdef VERILATOR
	DifftestInstrCommit DifftestInstrCommit(
		.clock              (clk),
		.coreid             (csr_regfile.mhartid[7:0]),
		.index              (0),
		.valid              (handin),
		.pc                 (dataW.pc),
		.instr              (0),
		.skip               (dataW.ctl.memwrite & ~dataW.mem_addr[31]),
		.isRVC              (0),
		.scFailed           (0),
		.wen                (dataW.ctl.regwrite),
		.wdest              ({3'b0, dataW.dst}),
		.wdata              (dataW.result)
	);
	      
	DifftestArchIntRegState DifftestArchIntRegState (
		.clock              (clk),
		.coreid             (csr_regfile.mhartid[7:0]),
		.gpr_0              (regfile.regs_nxt[0]),
		.gpr_1              (regfile.regs_nxt[1]),
		.gpr_2              (regfile.regs_nxt[2]),
		.gpr_3              (regfile.regs_nxt[3]),
		.gpr_4              (regfile.regs_nxt[4]),
		.gpr_5              (regfile.regs_nxt[5]),
		.gpr_6              (regfile.regs_nxt[6]),
		.gpr_7              (regfile.regs_nxt[7]),
		.gpr_8              (regfile.regs_nxt[8]),
		.gpr_9              (regfile.regs_nxt[9]),
		.gpr_10             (regfile.regs_nxt[10]),
		.gpr_11             (regfile.regs_nxt[11]),
		.gpr_12             (regfile.regs_nxt[12]),
		.gpr_13             (regfile.regs_nxt[13]),
		.gpr_14             (regfile.regs_nxt[14]),
		.gpr_15             (regfile.regs_nxt[15]),
		.gpr_16             (regfile.regs_nxt[16]),
		.gpr_17             (regfile.regs_nxt[17]),
		.gpr_18             (regfile.regs_nxt[18]),
		.gpr_19             (regfile.regs_nxt[19]),
		.gpr_20             (regfile.regs_nxt[20]),
		.gpr_21             (regfile.regs_nxt[21]),
		.gpr_22             (regfile.regs_nxt[22]),
		.gpr_23             (regfile.regs_nxt[23]),
		.gpr_24             (regfile.regs_nxt[24]),
		.gpr_25             (regfile.regs_nxt[25]),
		.gpr_26             (regfile.regs_nxt[26]),
		.gpr_27             (regfile.regs_nxt[27]),
		.gpr_28             (regfile.regs_nxt[28]),
		.gpr_29             (regfile.regs_nxt[29]),
		.gpr_30             (regfile.regs_nxt[30]),
		.gpr_31             (regfile.regs_nxt[31])
	);

    DifftestTrapEvent DifftestTrapEvent(
		.clock              (clk),
		.coreid             (csr_regfile.mhartid[7:0]),
		.valid              (0),
		.code               (0),
		.pc                 (0),
		.cycleCnt           (0),
		.instrCnt           (0)
	);

	DifftestCSRState DifftestCSRState(
		.clock              (clk),
		.coreid             (csr_regfile.mhartid[7:0]),
		.priviledgeMode     (privilege_mode_nxt),
		.mstatus            (csr_regfile.mstatus_nxt & MSTATUS_MASK),
		.sstatus            (csr_regfile.sstatus_nxt & SSTATUS_MASK),
		.mepc               (csr_regfile.mepc_nxt),
		.sepc               (0),
		.mtval              (csr_regfile.mtval_nxt),
		.stval              (0),
		.mtvec              (csr_regfile.mtvec_nxt & MTVEC_MASK),
		.stvec              (0),
		.mcause             (csr_regfile.mcause_nxt),
		.scause             (0),
		.satp               (csr_regfile.satp_nxt),
		.mip                (csr_regfile.mip_nxt & MIP_MASK),
		.mie                (csr_regfile.mie_nxt),
		.mscratch           (csr_regfile.mscratch_nxt),
		.sscratch           (0),
		.mideleg            (0),
		.medeleg            (0)
	);
`endif
endmodule
`endif
